module CPU
  (
   input  clk,
   input  inM [15:0],
   input  instruction [15:0],
   input  reset,
   output outM [15:0],
   output writeM,
   output addressM [15:0],
   output pc [15:0]
   );

   // TODO

endmodule // CPU


module ALU_tb();
   reg [15:0]  x;
   reg [15:0]  y;
   reg 	 zx;
   reg 	 nx;
   reg 	 zy;
   reg 	 ny;
   reg 	 f;
   reg 	 no;
   wire [15:0] out;
   wire 	 zr;
   wire 	 ng;

endmodule // ALU_tb

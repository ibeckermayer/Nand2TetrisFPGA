module CPU
  (
   input 	 clk,
   input [15:0]  inM,
   input [15:0]  instruction,
   input 	 reset,
   output [15:0] outM,
   output 	 writeM,
   output [15:0] addressM,
   output [15:0] pc
   );

   // TODO

endmodule // CPU

